module option_parser

const (
	helper_short = '-h'
	helper_long  = "--help"
	align_left   = 4
	align_middle = 33
)
