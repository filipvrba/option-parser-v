module option_parser

type Callback = fn (string)
